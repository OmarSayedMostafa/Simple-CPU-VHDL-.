----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:33:05 05/04/2016 
-- Design Name: 
-- Module Name:    FullAdder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FullAdder is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Carry : in  STD_LOGIC;
           OCarry : out  STD_LOGIC;
           O : out  STD_LOGIC);
end FullAdder;

architecture Behavioral of FullAdder is
signal tmp: std_logic_vector ( 1 downto 0 );
begin
 tmp <= ( '0' & A ) + ( '0' & B ) + ( '0' & Carry );

  O <= tmp(0);
  OCarry <= tmp(1);


end Behavioral;

